library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity wb_slave_arbiter is
  port (
	 -- Master to slave signals
	 i_wb_cyc			: in	std_logic;
	 i_wb_stb			: in	std_logic;
	 i_wb_we			: in	std_logic;
	 i_wb_addr			: in	std_logic_vector(31 downto 0);
	 i_wb_data			: in	std_logic_vector(31 downto 0);
	 i_wb_sel			: in	std_logic_vector( 3 downto 0);
	 o_wb_stall			: out std_logic;
	 o_wb_ack			: out std_logic;
	 o_wb_data			: out std_logic_vector(31 downto 0);
	 -- BRAM
	 o_wb_bram_cyc		: out std_logic;
	 o_wb_bram_stb		: out std_logic;
	 o_wb_bram_we		: out std_logic;
	 o_wb_bram_addr		: out std_logic_vector(31 downto 0);
	 o_wb_bram_data		: out std_logic_vector(31 downto 0);
	 o_wb_bram_sel		: out std_logic_vector( 3 downto 0);
	 i_wb_bram_stall	: in  std_logic;
	 i_wb_bram_ack		: in  std_logic;
	 i_wb_bram_data		: in  std_logic_vector(31 downto 0);
	 -- SDRAM
	 o_wb_sdram_cyc		: out std_logic;
	 o_wb_sdram_stb		: out std_logic;
	 o_wb_sdram_we		: out std_logic;
	 o_wb_sdram_addr	: out std_logic_vector(20 downto 0);
	 o_wb_sdram_data	: out std_logic_vector(31 downto 0);
	 o_wb_sdram_sel		: out std_logic_vector( 3 downto 0);
	 i_wb_sdram_stall	: in  std_logic;
	 i_wb_sdram_ack		: in  std_logic;
	 i_wb_sdram_data	: in  std_logic_vector(31 downto 0);
	 -- MMAP
	 o_wb_mmap_cyc		: out std_logic;
	 o_wb_mmap_stb		: out std_logic;
	 o_wb_mmap_we		: out std_logic;
	 o_wb_mmap_addr	: out std_logic_vector(31 downto 0);
	 o_wb_mmap_data	: out std_logic_vector(31 downto 0);
	 o_wb_mmap_sel		: out std_logic_vector( 3 downto 0);
	 i_wb_mmap_stall	: in  std_logic;
	 i_wb_mmap_ack		: in  std_logic;
	 i_wb_mmap_data	: in  std_logic_vector(31 downto 0);
	 -- ROM
	 o_wb_brom_cyc		: out std_logic;
	 o_wb_brom_stb		: out std_logic;
	 o_wb_brom_we		: out std_logic;
	 o_wb_brom_addr	: out std_logic_vector(31 downto 0);
	 o_wb_brom_data	: out std_logic_vector(31 downto 0);
	 o_wb_brom_sel		: out std_logic_vector( 3 downto 0);
	 i_wb_brom_stall	: in  std_logic;
	 i_wb_brom_ack		: in  std_logic;
	 i_wb_brom_data	: in  std_logic_vector(31 downto 0)
    );
end entity;

architecture rtl of wb_slave_arbiter is
	
	type t_slave is (BROM, BRAM, SDRAM, MMAP, SEGFAULT);
	signal s_slave : t_slave;
	
begin

	-- BROM			0x000000 - 0x000FFF ( 4KiB)
	-- BRAM			0x001000 - 0x00BFFF (20KiB)
	-- Peripherals	0x008000 - 0x00BFFF (16KiB)
	-- SDRAM 		0x00C000 - 0x10BFFF ( 1MiB)

	s_slave <= BROM when i_wb_addr < 16#1000# else
				  BRAM when i_wb_addr < 16#8000# else
				  MMAP when i_wb_addr < 16#C000# else
				  SDRAM when i_wb_addr < 16#10C000# else
				  SEGFAULT;

	-- Slave to Master outputs
	o_wb_stall <= i_wb_brom_stall when s_slave = BROM else
					  i_wb_bram_stall when s_slave = BRAM else
					  i_wb_mmap_stall when s_slave = MMAP else
					  i_wb_sdram_stall when s_slave = SDRAM else
					  '0';
	o_wb_ack <= i_wb_brom_ack when s_slave = BROM else
					i_wb_bram_ack when s_slave = BRAM else
					i_wb_mmap_ack when s_slave = MMAP else
					i_wb_sdram_ack when s_slave = SDRAM else
					'0';
	o_wb_data <= i_wb_brom_data when s_slave = BROM else
					 i_wb_bram_data when s_slave = BRAM else
					 i_wb_mmap_data when s_slave = MMAP else
					 i_wb_sdram_data when s_slave = SDRAM else
					 (others => '0');
	
	-- BROM
	o_wb_brom_cyc <= i_wb_cyc when s_slave = BROM else '0';
	o_wb_brom_stb <= i_wb_stb when s_slave = BROM else '0';
	o_wb_brom_we <= i_wb_we when s_slave = BROM else '0';
	o_wb_brom_addr <= i_wb_addr when s_slave = BROM else (others => '0');
	o_wb_brom_data <= i_wb_data when s_slave = BROM else (others => '0');
	o_wb_brom_sel <= i_wb_sel when s_slave = BROM else (others => '0');
    
	-- BRAM
	o_wb_bram_cyc <= i_wb_cyc when s_slave = BRAM else '0';
	o_wb_bram_stb <= i_wb_stb when s_slave = BRAM else '0';
	o_wb_bram_we <= i_wb_we when s_slave = BRAM else '0';
	o_wb_bram_addr <= i_wb_addr - 16#1000# when s_slave = BRAM else (others => '0');
	o_wb_bram_data <= i_wb_data when s_slave = BRAM else (others => '0');
	o_wb_bram_sel <= i_wb_sel when s_slave = BRAM else (others => '0');

	-- MMAP Peripherals
	o_wb_mmap_cyc <= i_wb_cyc when s_slave = MMAP else '0';
	o_wb_mmap_stb <= i_wb_stb when s_slave = MMAP else '0';
	o_wb_mmap_we <= i_wb_we when s_slave = MMAP else '0';
	o_wb_mmap_addr <= i_wb_addr - 16#8000# when s_slave = MMAP else (others => '0');
	o_wb_mmap_data <= i_wb_data when s_slave = MMAP else (others => '0');
	o_wb_mmap_sel <= i_wb_sel when s_slave = MMAP else (others => '0');

	-- SDRAM
	o_wb_sdram_cyc <= i_wb_cyc when s_slave = SDRAM else '0';
	o_wb_sdram_stb <= i_wb_stb when s_slave = SDRAM else '0';
	o_wb_sdram_we <= i_wb_we when s_slave = SDRAM else '0';
	o_wb_sdram_addr <= i_wb_addr(20 downto 0) when s_slave = SDRAM else (others => '0');
	o_wb_sdram_data <= i_wb_data when s_slave = SDRAM else (others => '0');
	o_wb_sdram_sel <= i_wb_sel when s_slave = SDRAM else (others => '0');

end architecture;
